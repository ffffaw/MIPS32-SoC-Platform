module UART_RX (
	input wire clk,
	input wire rstn,
	input wire b_tick,        // Baud generator tick
	input wire rx,            // RS-232 data port
	
	output reg rx_done,       // transfer completed
	output wire [7:0] dout,   // output data

	input parity_check// ================================================================
);

	// STATE DEFINES  
	localparam [1:0] idle_st = 2'b00;
	localparam [1:0] start_st = 2'b01;
	localparam [1:0] data_st = 2'b11;
	localparam [1:0] stop_st = 2'b10;

	// Internal Signals  
	reg [1:0] current_state;
	reg [1:0] next_state;
	reg [3:0] b_reg;// baud-rate/over sampling counter
	reg [3:0] b_next;
	reg [2:0] count_reg;// data-bit counter
	reg [2:0] count_next;
	reg [7:0] data_reg;// data register
	reg [7:0] data_next;
	
	// State Machine  
	always @(posedge clk, negedge rstn)
	begin
		if(!rstn)
		begin
			current_state <= idle_st;
			b_reg <= 0;
			count_reg <= 0;
			data_reg <=0;
		end
		else
		begin
			current_state <= next_state;
			b_reg <= b_next;
			count_reg <= count_next;
			data_reg <= data_next;
		end
	end

	// Next State Logic 
	always @(*)
	begin
		next_state = current_state;
		b_next = b_reg;
		count_next = count_reg;
		data_next = data_reg;
		rx_done = 1'b0;

		case(current_state)
		idle_st:
			if(~rx)
			begin
				next_state = start_st;
				b_next = 0;
			end
			
		start_st:
			if(b_tick)
				if(b_reg == 3)
					begin
						next_state = data_st;
						b_next = 0;
						count_next = 0;
					end
				else
					b_next = b_reg + 1'b1;
				
		data_st:
			if(b_tick)
				if(b_reg == 3)
				begin
					b_next = 0;
					data_next = {rx, data_reg[7:1]};
					if(count_next == 7) // 8 Data bits
						next_state = stop_st;
					else
						count_next = count_reg + 1'b1;
				end
			else
				b_next = b_reg + 1;
				
		stop_st:
			if(b_tick)
				if(b_reg == 3) // One stop bit
					begin
						next_state = idle_st;
						// rx_done = 1'b1;
						// ================================================================ parity check below
						if(parity_check == 0)
						begin
							rx_done = 1'b1;
						end
						else
						begin
							if((data_reg[7] ^ data_reg[6] ^ data_reg[5] ^ data_reg[4] ^ data_reg[3] ^
								data_reg[2] ^ data_reg[1] ^ data_reg[0]) == 1)
							begin
								rx_done = 1'b1;
							end
							else
							begin
								rx_done = 1'b0;
							end
						end
						// ================================================================ parity check above
						
					end
				else
				b_next = b_reg + 1;
		endcase
	end
	
	assign dout = data_reg;
	
endmodule


